LIBRARY IEEE;

package constants is
    constant BITS_ARCH   : integer ;
    constant SEL_ARCH    : integer := 4;
    constant SEG7_AMOUNT : integer := 2;
end constants;
